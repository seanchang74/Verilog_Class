module matrix2 (clk,reset,segout,scanout);

input clk,reset;
output reg[7:0] segout;
output reg[2:0] scanout;

reg[25:0] cnt_scan;//
reg[6:0] i=0;

reg clk1;
reg [7:0] q[0:7] ;

//------------------ clock running -----------------------
always@(posedge clk or negedge reset)
begin
	if(!reset) begin
		cnt_scan<=0;
	end
	else begin
		cnt_scan<=cnt_scan+1;
		if (cnt_scan == 6250000) begin
			cnt_scan <=0;
			clk1 = ~clk1;
		end
	end
end

//---------modify display digit ----------
always @(posedge clk1 , negedge reset)
begin

	if (reset == 0)
	begin
		q[0] = 8'b11111111;
		q[1] = 8'b11111111;
		q[2] = 8'b11111111;
		q[3] = 8'b11111111;
		q[4] = 8'b11111111;
		q[5] = 8'b11111111;
		q[6] = 8'b11111111;
		q[7] = 8'b11111111;				
	end
	else begin
		case(i)
		1:
		begin
		q[0] <= 8'b11101111;
		i = i + 1;
		end
		2:
		begin
		q[0] <= 8'b11011111;
		q[1] <= 8'b11011111;
		i = i + 1;
		end
		3:
		begin
		q[0] <= 8'b10111111;
		q[1] <= 8'b10111111;
		q[2] <= 8'b10111111;
		i = i+1;
		end
		4:
		begin
		q[0] <= 8'b01111111;
		q[1] <= 8'b01111111;
		q[2] <= 8'b01111111;
		q[3] <= 8'b01111111;
		i = i+1;
		end
		5:
		begin
		q[0] <= 8'b11111111;
		q[1] <= 8'b01111111;
		q[2] <= 8'b01111111;
		q[3] <= 8'b01111111;
		q[4] <= 8'b01111111;
		i = i+1;
		end
		6:
		begin
		q[1] <= 8'b11111111;
		q[2] <= 8'b01111111;
		q[3] <= 8'b01111111;
		q[4] <= 8'b01111111;
		q[5] <= 8'b01111111;
		i = i+1;
		end
		7:
		begin
		q[2] <= 8'b11111111;
		q[3] <= 8'b01111111;
		q[4] <= 8'b01111111;
		q[5] <= 8'b01111111;
		q[6] <= 8'b01111111;
		i = i+1;
		end
		8:
		begin
		q[3] <= 8'b11111111;
		q[4] <= 8'b01111111;
		q[5] <= 8'b01111111;
		q[6] <= 8'b01111111;
		q[7] <= 8'b01111111;
		i = i+1;
		end
		9:
		begin
		q[0] <= 8'b11101111;
		i = i+1;
		end
		10:
		begin
		q[0] <= 8'b11100111;
		q[1] <= 8'b11101111;
		i = i+1;
		end
		11:
		begin
		q[0] <= 8'b11101111;
		q[1] <= 8'b11100111;
		q[2] <= 8'b11101111;
		i = i+1;
		end
		12:
		begin
		q[0] <= 8'b11011111;
		q[1] <= 8'b10001111;
		q[2] <= 8'b11111111;
		i = i+1;
		end
		13:
		begin
		q[0] <= 8'b11111111;
		q[1] <= 8'b11011111;
		q[2] <= 8'b10001111;
		i = i+1;
		end
		14:
		begin
		q[1] <= 8'b11111111;
		q[2] <= 8'b11011111;
		q[3] <= 8'b10001111;
		i = i+1;
		end
		15:
		begin
		q[2] <= 8'b11111111;
		q[3] <= 8'b11011111;
		q[4] <= 8'b00001111;
		i = i+1;
		end
		16:
		begin
		q[3] <= 8'b11111111;
		q[4] <= 8'b01011111;
		q[5] <= 8'b00001111;
		i = i+1;
		end
		17:
		begin
		q[4] <= 8'b01111111;
		q[5] <= 8'b01011111;
		q[6] <= 8'b00001111;
		i = i+1;
		end
		18:
		begin
		q[5] <= 8'b01111111;
		q[6] <= 8'b01011111;
		q[7] <= 8'b00001111;
		i = i+1;
		end
		19:
		begin
		q[0] <= 8'b11101111;
		i = i+1;
		end
		20:
		begin
		q[0] <= 8'b11101111;
		q[1] <= 8'b11101111;
		i = i+1;
		end
		21:
		begin
		q[0] <= 8'b11100111;
		q[1] <= 8'b11110111;
		q[2] <= 8'b11110111;
		i = i+1;
		end
		22:
		begin
		q[0] <= 8'b11111011;
		q[1] <= 8'b11100011;
		q[2] <= 8'b11111111;
		i = i+1;
		end
		23:
		begin
		q[0] <= 8'b11111111;
		q[1] <= 8'b11111101;
		q[2] <= 8'b11110001;
		i = i+1;
		end
		24:
		begin
		q[1] <= 8'b11111111;
		q[2] <= 8'b11111110;
		q[3] <= 8'b11111000;
		i = i+1;
		end
		25:
		begin
		q[2] <= 8'b11111111;
		q[3] <= 8'b11111110;
		q[4] <= 8'b01111000;
		i = i+1;
		end
		26:
		begin
		q[3] <= 8'b11111111;
		q[4] <= 8'b01111110;
		q[5] <= 8'b01111000;
		i = i+1;
		end
		27:
		begin
		q[4] <= 8'b01111111;
		q[5] <= 8'b01111110;
		q[6] <= 8'b01011000;
		i = i+1;
		end
		28:
		begin
		q[5] <= 8'b01111111;
		q[6] <= 8'b01011110;
		q[7] <= 8'b00001000;
		i = i+1;
		end
		29:
		begin
		q[0] <= 8'b11101111;
		i = i+1;
		end
		30:
		begin
		q[0] <= 8'b11100111;
		q[1] <= 8'b11101111;
		i = i+1;
		end
		31:
		begin
		q[0] <= 8'b11101111;
		q[1] <= 8'b11100111;
		q[2] <= 8'b11101111;
		i = i+1;
		end
		32:
		begin
		q[0] <= 8'b11111111;
		q[1] <= 8'b11110111;
		q[2] <= 8'b11110011;
		q[3] <= 8'b11110111;
		i = i+1;
		end
		33:
		begin
		q[1] <= 8'b11111111;
		q[2] <= 8'b11110111;
		q[3] <= 8'b11110011;
		q[4] <= 8'b01110111;
		i = i+1;
		end
		34:
		begin
		q[2] <= 8'b11111111;
		q[3] <= 8'b11110111;
		q[4] <= 8'b01110011;
		q[5] <= 8'b01110111;
		i = i+1;
		end
		35:
		begin
		q[3] <= 8'b11111111;
		q[4] <= 8'b01110111;
		q[5] <= 8'b01110011;
		q[6] <= 8'b01010110;
		i = i+1;
		end
		36:
		begin
		q[4] <= 8'b01111111;
		q[5] <= 8'b01110111;
		q[6] <= 8'b01010010;
		q[7] <= 8'b00000000;
		i = i+1;
		end
		37:
		begin
		q[4] <= 8'b01111111;
		q[5] <= 8'b01110111;
		q[6] <= 8'b01010010;
		q[7] <= 8'b11111111;
		i = i+1;
		end
		38:
		begin
		q[4] <= 8'b11111111;
		q[5] <= 8'b01111111;
		q[6] <= 8'b01110111;
		q[7] <= 8'b01010010;		
		i = i+1;
		end
		39:
		begin
		q[0] <= 8'b11101111;
		i = i+1;
		end
		40:
		begin
		q[0] <= 8'b11101111;
		q[1] <= 8'b11101111;
		i = i+1;
		end
		41:
		begin
		q[0] <= 8'b11001111;
		q[1] <= 8'b11011111;
		q[2] <= 8'b11011111;
		i = i+1;
		end
		42:
		begin
		q[0] <= 8'b11111111;
		q[1] <= 8'b11001111;
		q[2] <= 8'b11011111;
		q[3] <= 8'b11011111;
		i = i+1;
		end
		43:
		begin
		q[1] <= 8'b11111111;
		q[2] <= 8'b10011111;
		q[3] <= 8'b10111111;
		q[4] <= 8'b10111111;
		i = i+1;
		end
		44:
		begin
		q[2] <= 8'b11111111;
		q[3] <= 8'b10011111;
		q[4] <= 8'b10111111;
		q[5] <= 8'b00111111;
		i = i+1;
		end
		45:
		begin
		q[3] <= 8'b11111111;
		q[4] <= 8'b10011111;
		q[5] <= 8'b00111111;
		q[6] <= 8'b00110111;
		i = i+1;
		end
		46:
		begin
		q[4] <= 8'b11111111;
		q[5] <= 8'b00011111;
		q[6] <= 8'b00110111;
		q[7] <= 8'b00010010;
		i = i+1;
		end
		47:
		begin
		q[0] <= 8'b11101111;
		i = i+1;
		end
		48:
		begin
		q[0] <= 8'b11001111;
		q[1] <= 8'b11101111;
		i = i+1;
		end
		49:
		begin
		q[0] <= 8'b11101111;
		q[1] <= 8'b11100111;
		q[2] <= 8'b11110111;
		i = i+1;
		end
		50:
		begin
		q[0] <= 8'b11111111;
		q[1] <= 8'b11110111;
		q[2] <= 8'b11110011;
		q[3] <= 8'b11111011;
		i = i+1;
		end
		51:
		begin
		q[1] <= 8'b11111111;
		q[2] <= 8'b11111011;
		q[3] <= 8'b11111001;
		q[4] <= 8'b11111101;
		i = i+1;
		end
		52:
		begin
		q[2] <= 8'b11111111;
		q[3] <= 8'b11111011;
		q[4] <= 8'b11111001;
		q[5] <= 8'b00011101;
		i = i+1;
		end
		53:
		begin
		q[3] <= 8'b11111111;
		q[4] <= 8'b11111011;
		q[5] <= 8'b00011001;
		q[6] <= 8'b00110101;
		i = i+1;
		end
		54:
		begin
		q[4] <= 8'b11111111;
		q[5] <= 8'b00011011;
		q[6] <= 8'b00110001;
		q[7] <= 8'b00010000;
		i = i+1;
		end
		55:
		begin
		q[0] <= 8'b10000111;
		i = i+1;
		end
		56:
		begin
		q[0] <= 8'b11101111;
		q[1] <= 8'b11101111;
		i = i+1;
		end
		57:
		begin
		q[0] <= 8'b11101111;
		q[1] <= 8'b11101111;
		q[2] <= 8'b11101111;
		i = i+1;
		end
		58:
		begin
		q[0] <= 8'b11101111;
		q[1] <= 8'b11101111;
		q[2] <= 8'b11101111;
		q[3] <= 8'b11101111;
		i = i+1;
		end
		59:
		begin
		q[0] <= 8'b11111111;
		q[1] <= 8'b11101111;
		q[2] <= 8'b11101111;
		q[3] <= 8'b11101111;
		q[4] <= 8'b11101111;
		i = i+1;
		end
		60:
		begin
		q[1] <= 8'b11111111;
		q[2] <= 8'b11101111;
		q[3] <= 8'b11101111;
		q[4] <= 8'b11101111;
		q[5] <= 8'b00001011;
		i = i+1;
		end
		61:
		begin
		q[2] <= 8'b11111111;
		q[3] <= 8'b11101111;
		q[4] <= 8'b11101111;
		q[5] <= 8'b00001011;
		q[6] <= 8'b00100001;
		i = i+1;
		end
		62:
		begin
		q[3] <= 8'b11111111;
		q[4] <= 8'b11101111;
		q[5] <= 8'b00001011;
		q[6] <= 8'b00100001;
		q[7] <= 8'b00000000;
		i = i+1;
		end
		63:
		begin
		q[7] <= 8'b11111111;
		i = i+1;
		end
		64:
		begin
		q[4] <= 8'b11111111;
		q[5] <= 8'b11101111;
		q[6] <= 8'b00001011;
		q[7] <= 8'b00100001;
		i = i+1;
		end
		65:
		begin
		q[4] <= 8'b11111111;
		q[5] <= 8'b11101111;
		q[6] <= 8'b00001011;
		q[7] <= 8'b00100001;
		i = i+1;
		end
		default:
		begin
		q[0] <= 8'b11111111;
		q[1] <= 8'b11111111;
		q[2] <= 8'b11111111;
		q[3] <= 8'b11111111;
		q[4] <= 8'b11111111;
		q[5] <= 8'b11111111;
		q[6] <= 8'b11111111;
		q[7] <= 8'b11111111;
		i = 1;	
		end		
		endcase
	end
end
//-----------scan and display 7-SEG-------------
always@(cnt_scan[15:13])
begin
	scanout <= cnt_scan[15:13];
end

	always@(scanout) //
	begin
		case(scanout)
			0: segout=q[0];
			1: segout=q[1];
			2: segout=q[2];
			3: segout=q[3];
			4: segout=q[4];
			5: segout=q[5];
			6: segout=q[6];
			7: segout=q[7];
		default:
			segout=8'b11111111;
		endcase
	end

endmodule
